library IEEE;
use IEEE.std_logic_1164.all;

entity t_ff is
    port (
        
    );
end entity t_ff;